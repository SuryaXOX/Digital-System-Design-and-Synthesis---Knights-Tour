module cmd_proc_tb();

/* GLOBAL SIGNALS */
parameter FAST_SIM = 1;
// remote_comm
logic clk, rst_n;
logic [15:0] cmd;
logic send_cmd, resp_rdy, cmd_sent;
logic [7:0] resp;
// uart_wrapper
logic trmt;
logic tx_done;
// cmd_proc
logic lftIR, rghtIR, cntrIR;
logic fanfare_go, tour_go;
logic moving, rdy;
logic [9:0] frwrd;
logic [11:0] error;

/* INTERMEDIATE SIGNALS */
logic TX_RX, RX_TX;                     // remote-wrapper
logic INT, SS_n, SCLK, MOSI, MISO;      // spi-integrator
// integrator-cmd_proc
logic [11:0] heading;
logic heading_rdy;
logic strt_cal, cal_done;
// wrapper-cmd_proc
logic [15:0] cmd_wrapper;
logic cmd_rdy, clr_cmd_rdy;
logic send_resp;


/* INITIALIZING MODULES */
RemoteComm REMOTE_COMM(.clk(clk), .rst_n(rst_n), .RX(RX_TX), .TX(TX_RX), .cmd(cmd), .send_cmd(send_cmd), .cmd_sent(cmd_sent), .resp_rdy(resp_rdy), .resp(resp));
UART_wrapper WRAPPER(.clk(clk), .rst_n(rst_n), .clr_cmd_rdy(clr_cmd_rdy), .cmd_rdy(cmd_rdy), .cmd(cmd_wrapper), .trmt(send_resp), .resp(8'hA5), .tx_done(tx_done), .RX(TX_RX), .TX(RX_TX));
SPI_iNEMO3 SPI_NEMO(.SS_n(SS_n), .SCLK(SCLK), .MISO(MISO), .MOSI(MOSI), .INT(INT));
inert_intf INTEGRATOR(.clk(clk), .rst_n(rst_n), .lftIR(lftIR), .rghtIR(rghtIR), .moving(moving), .heading(heading), .strt_cal(strt_cal), .cal_done(cal_done), .rdy(heading_rdy), 
     .SS_n(SS_n), .SCLK(SCLK), .MISO(MISO), .MOSI(MOSI), .INT(INT));
cmd_proc #(FAST_SIM) CMD_PROC(.clk(clk), .rst_n(rst_n), .cmd(cmd_wrapper), .cmd_rdy(cmd_rdy), .clr_cmd_rdy(clr_cmd_rdy), .send_resp(send_resp), .strt_cal(strt_cal),
                .cal_done(cal_done), .heading(heading), .heading_rdy(heading_rdy), .lftIR(lftIR), .cntrIR(cntrIR), .rghtIR(rghtIR), .error(error),
				.frwrd(frwrd), .moving(moving), .tour_go(tour_go), .fanfare_go(fanfare_go));

initial begin
    // initializing signals
    clk = 1'b0;
    rst_n = 1'b0;
    send_cmd = 1'b0;
    cmd = 16'h0000;
    lftIR = 1'b0;
    rghtIR = 1'b0;
    trmt = 1'b0;
    cmd_rdy = 1'b0;

    @(posedge clk);
    @(negedge clk) rst_n = 1'b1;
    send_cmd = 1;
    @(posedge clk);
    @(negedge clk);
    send_cmd = 0;
   /* // asserting snd_cmd for one clock cycle
    @(posedge clk);
    strt_cal = 1'b1;
    @(posedge clk);
    strt_cal = 1'b0;
   */
    // waiting for cal_done and resp_rdy signals to be asserted
    fork
        // timeout
        begin: timeout1
            repeat(1000000) @(posedge clk);
            $display("ERROR: timed out waiting for cal_done to assert");
            $stop();
        end
        // watiting for cal_done
        begin
            @(posedge cal_done);
            disable timeout1;
        end
        // timeout
        begin: timeout2
            // wait
            repeat(1000000) @(posedge clk);
            $display("ERROR: timed out waiting for resp_rdy to assert");
            $stop();
        end
        // waiting for resp_rdy
        begin
            @(posedge resp_rdy);
            disable timeout2;
        end
    join
    
    $display("SUCCESS: got cal_done and resp_rdy asserted!");
    
    // SENDING NORTH CMD, 1
    @(posedge clk);
    cmd = 16'h2001;
    send_cmd = 1;
    @(posedge clk);
    @(negedge clk);
    send_cmd = 0;
   

    // waiting for cmd_sent
    fork
        begin: timeout3
            // wait
            repeat(100000) @(posedge clk);
            $display("ERROR: timed out waiting for cmd_sent to assert");
            $stop();
        end
        // waiting for cmd_sent
        begin
            @(posedge cmd_sent);
            //if(cmd_sent)
            disable timeout3;
        end
    join

    $display("SUCCESS: cmd_sent asserted!");
    
    // checking if frwrd is set properly
    if (frwrd!==10'h000) begin
        $display("frwrd should be 10'h000 but you got %h", frwrd);
        $stop();
    end
    
    $display("SUCCESS: frwrd is set properly!");

    // checking if frwrd increments properly
    repeat(10) @(posedge heading_rdy);
    if (frwrd !== (10'h120) && frwrd !== (10'h140)) begin
        $display("frwrd should be 10'h120 or 10'h140 but you got %h", frwrd);
        $stop();
    end
    
    $display("SUCCESS: frwrd is set properly to x120 or x140!");

    // making sure that moving signal is asserted
    if (!moving) begin
        $display("moving should be asserted but it is %h", moving);
        $stop();
    end

    // checking if frwrd is saturated
    repeat(20) @(posedge heading_rdy);
    if (~&frwrd[9:8]) begin
        $display("frwrd after few cycles should be maxed out but you got %h", frwrd);
        $stop();
    end

    // check if frwrd is still saturated after 'crossing one line', it should be saturated
    cntrIR = 1'b1;
    @(posedge clk);
    cntrIR = 1'b0;
    repeat(5) @(posedge clk);
    if (~&frwrd[9:8]) begin
        $display("frwrd after crossing 1 line should be maxed out but you got %h", frwrd);
        $stop();
    end

    // check if frwrd is still saturated after 'crossing second line', it should NOT be saturated
    cntrIR = 1'b1;
    @(posedge clk);         // NOT SURE HOW LONG THE PULSE SHOULD BE, DOUBLE CHECK
    cntrIR = 1'b0;
    repeat(5) @(posedge clk);
    if (&frwrd[9:8]) begin
        $display("frwrd after crossing 2 lines should not be maxed out but it is, you got %h", frwrd);
        $stop();
    end

    $display("SUCCESS: crossed 2 lines");

    // checking for resp_rdy
    fork
        begin: timeout4
            // wait
            repeat(100000) @(negedge clk);
            $display("ERROR: timed out waiting for resp_rdy to assert");
            $stop();
        end
        // waiting for resp_rdy
        begin
            @(posedge resp_rdy);
            disable timeout4;
        end
        // checking if frwrd reaches zero
        @(negedge |frwrd) $display("frwrd reached 0!");        
    join


    /* END OF MINIMUM TESTS */

    // rghtIR/lftIR test, SENDING NORTH CMD, 2
    
    cmd = 16'h2001;
    @(posedge clk);
    send_cmd = 1;
    @(posedge clk);
    @(negedge clk);
    send_cmd = 0;

    // waiting for cmd_sent
    fork
        begin: timeout5
            // wait
            repeat(100000) @(negedge clk);
            $display("ERROR: timed out waiting for cmd_sent to assert");
            $stop();
        end
        // waiting for cmd_sent
        begin
            @(posedge cmd_sent);
            disable timeout5;
        end
    join

    // checking if frwrd is set properly
    if (frwrd!==10'h000) begin
        $display("frwrd should be 10'h000 but you got %h", frwrd);
        $stop();
    end

    // checking if frwrd increments properly
    repeat(10) @(posedge heading_rdy);
    if (frwrd!==10'h120 && frwrd!==10'h140) begin
        $display("frwrd should be 10'h120 or 10'h140 but you got %h", frwrd);
        $stop();
    end

    // making sure that moving signal is asserted
    if (!moving) begin
        $display("moving should be asserted but it is %h", moving);
        $stop();
    end

    // checking if frwrd is saturated
    repeat(20) @(posedge heading_rdy);
    if (~&frwrd[9:8]) begin
        $display("frwrd after few cycles should be maxed out but you got %h", frwrd);
        $stop();
    end

    // sending lftIR pulse, recording error value before that

    rghtIR = 1'b1;
    repeat(600000) @(posedge clk);
    rghtIR = 1'b0;

    // checking for disturbance in error by looking at wave difference
    // TODO: make self-checking

    $stop();
end

always
    #5 clk = ~clk;

endmodule





